/*
 * The SPI is used as an interface between the SOM and
 * the FPGA in order to (from the point of view of the FPGA):
 *   - Receive a new configuration for the drivers
 *   - Transmit rotation information given by the Hall effect
 *   sensors to the SBC
 */

module spi_decoder (
    input  nrst,
    input  clk,

    input  valid,
    input  [391:0] data_mosi,
    input  [10:0]  data_len_bytes,
    output [47:0] data_miso,

    // Data generated by the Hall sensor module
    input [15:0] rotation_data,
    input [15:0] speed_data,
    input [31:0] debug_data,
    output [47:0] configuration,

    output new_config_available,
    output rgb_enable,

    // Mux statuses
    output [7:0] mux,

    output [47:0] driver_data [29:0],
    output [431:0] debug_driver,
    output         debug_driver_override_lut,

    // Signals that the topmodule should use debugging data signals from the spi_decoder
    output manage
);

localparam CONFIG_COMMAND = 'hBF;
localparam ROTATION_COMMAND = 'h4C;
localparam SPEED_COMMAND = 'h4D;
localparam DISABLE_RGB_COMMAND = 'hD0;
localparam ENABLE_RGB_COMMAND = 'hE0;
localparam DEBUG_COMMAND = 'hDE;
localparam ENABLE_MUX_COMMAND = 'hE1;
localparam DISABLE_MUX_COMMAND = 'hD1;
localparam DRIVER_DATA_COMMAND = 'hDD;
localparam DRIVER_COMMAND_RGB = 'hEE;   // Still uses the LUTs
localparam DRIVER_COMMAND_POKER = 'hEF; // Overrides output LUTs
localparam MANAGE_COMMAND = 'hFA;
localparam RELEASE_COMMAND = 'hFE;

`include "drivers_conf.svh"

logic [391:0] last_cmd_read;
logic [10:0] last_cmd_len_bytes;
logic last_valid;

always_ff @(posedge clk or negedge nrst)
    if (~nrst) begin
        last_cmd_read <= '0;
        last_cmd_len_bytes <= '0;
        last_valid <= '0;
    end else begin
        last_valid <= valid;
        if(valid) begin
            last_cmd_read <= data_mosi;
            last_cmd_len_bytes <= data_len_bytes;
        end
    end

always_ff @(posedge clk or negedge nrst)
    if (~nrst) begin
        configuration <= serialized_conf;
        new_config_available <= 1;       // This will be high for one cycle (STALL)
        rgb_enable <= 0;
        mux <= '0;
        debug_driver <= '0;
        debug_driver_override_lut <= '0;
        manage <= '0;
        for (int i=0; i<30; ++i) begin
            driver_data[i] <= '0;
        end
    end else begin
        new_config_available <= '0;
        if (last_valid) begin
            if (last_cmd_len_bytes == 7 && last_cmd_read[55:48] == CONFIG_COMMAND) begin
                configuration <= last_cmd_read[47:0];
                new_config_available <= '1;
                data_miso <= configuration;
            end else if (last_cmd_len_bytes == 1
                         && last_cmd_read[7:0] == MANAGE_COMMAND) begin
                manage <= 1;
            end else if (last_cmd_len_bytes == 1
                         && last_cmd_read[7:0] == RELEASE_COMMAND) begin
                manage <= 0;
            end else if (last_cmd_len_bytes == 1
                         && last_cmd_read[7:0] == CONFIG_COMMAND) begin
                data_miso <= configuration;
            end else if (last_cmd_len_bytes == 1
                         && last_cmd_read[7:0] == ROTATION_COMMAND) begin
                data_miso[47:32] <= rotation_data;
            end else if (last_cmd_len_bytes == 1
                         && last_cmd_read[7:0] == SPEED_COMMAND) begin
                data_miso[47:32] <= speed_data;
            end else if (last_cmd_len_bytes == 1
                         && last_cmd_read[7:0] == DEBUG_COMMAND) begin
                data_miso <= {16'b0, debug_data};
            end else if (last_cmd_len_bytes == 49
                         && last_cmd_read[391:384] == DRIVER_COMMAND_RGB) begin
                debug_driver <= last_cmd_read[383:0];
                debug_driver_override_lut <= 0;
            end else if (last_cmd_len_bytes == 55
                         && last_cmd_read[439:432] == DRIVER_COMMAND_POKER) begin
                debug_driver <= last_cmd_read[431:0];
                debug_driver_override_lut <= 1;
            end else if (last_cmd_len_bytes == 1
                         && last_cmd_read[7:0] == ENABLE_RGB_COMMAND) begin
                rgb_enable <= '1;
            end else if (last_cmd_len_bytes == 1
                         && last_cmd_read[7:0] == DISABLE_RGB_COMMAND) begin
                rgb_enable <= '0;
            end else if (last_cmd_len_bytes == 2
                         && last_cmd_read[15:8] == ENABLE_MUX_COMMAND) begin
                mux[last_cmd_read[2:0]] <= 1;
            end else if (last_cmd_len_bytes == 2
                         && last_cmd_read[15:8] == DISABLE_MUX_COMMAND) begin
                mux[last_cmd_read[2:0]] <= 0;
            end else if (last_cmd_len_bytes == 8
                         && last_cmd_read[63:56] == DRIVER_DATA_COMMAND) begin
                if (last_cmd_read[55:48] < 8'd30)
                    driver_data[last_cmd_read[52:48]] <= last_cmd_read[47:0];
            end
        end
    end

endmodule
