/*
 * The SPI is used as an interface between the SOM and
 * the FPGA in order to (from the point of view of the FPGA):
 *   - Receive a new configuration for the drivers
 *   - Transmit rotation information given by the Hall effect
 *   sensors to the SBC
 */

module spi_slave(
    input  nrst,

    input  spi_clk,
    input  spi_ss,
    input  spi_mosi,
    output spi_miso,

    // Data generated by the Hall sensor module
    input [15:0] rotation_data,

    output [47:0] config_out,
    output new_config_available,
    output rgb_enable
);

localparam CONFIG_COMMAND = 191;
localparam ROTATION_COMMAND = 76;
localparam DISABLE_RGB_COMMAND = 'hD0;
localparam ENABLE_RGB_COMMAND = 'hE0;
localparam DEFAULT_CONFIG_DATA = 'hff;

/*
 * ReceiveRegister is a shift register for the received byte
 * TransmitRegister is a shift register for the byte to be transmitted
 */
logic [7:0] receive_register, transmit_register;

/*
 * shift_counter keeps trace of the number of times the receive_register is
 * shifted
 */
logic [3:0] shift_counter;

// Counter that counts the number of configuration bytes received
logic [2:0] config_byte_counter;

/*
 * State and counter for the transmission,
 */
enum logic [1:0] {NO_TRANSMISSION, FIRST_BYTE, SECOND_BYTE} transmission_step;

// 48-bit register that stores the received configuration
/* verilator lint_off UNUSED */
logic [47:0] configuration;
/* verilatro lint_off WIDTH */
assign config_out = configuration;

// Send bit of the transmission shift register when in transmission mode
assign spi_miso = transmission_step == NO_TRANSMISSION ? 1'b1 : transmit_register[7];

/*
 * Process for the receiving part:
 * The master sends data through spi_mosi while ss is low,
 * it is stored in the receive_register, which is then
 * shifted.
 */
always_ff @(posedge spi_clk or negedge nrst) begin
    if (~nrst) begin
        shift_counter <= '0;
    end else begin
        if (~spi_ss) begin
            // Shift the receive register
            receive_register[7:1] <= receive_register[6:0];
            // Store the incoming spi_mosi data in the receive register LSB
            receive_register[0] <= spi_mosi;
            shift_counter <= shift_counter + 1'b1;
            if (shift_counter == 7) begin
                shift_counter <= '0;
            end
        end else begin
            shift_counter <= '0;
        end
    end
end

/*
 * Process for the receiver logic.
 * It outputs the received bytes in the right order
 * in the output configuration.
 */
always_ff @(posedge spi_clk or negedge nrst) begin
    if (~nrst) begin
        config_byte_counter <= 0;
        new_config_available <= 0;
    end else begin
        if (config_byte_counter == 0 && shift_counter == 0) begin
            case (receive_register)
                CONFIG_COMMAND: begin
                    config_byte_counter <= 1;
                    configuration[7:0] <= receive_register;
                end
                DISABLE_RGB_COMMAND: begin
                    rgb_enable <= 0;
                end
                ENABLE_RGB_COMMAND: begin
                    rgb_enable <= 1;
                end
            endcase
        end
        if (config_byte_counter > 0 && shift_counter == 0) begin
            configuration[(config_byte_counter-1)*8 +: 8] <= receive_register;
            if (config_byte_counter == 6) begin
                /*
                * When the whole new configuration is received, reset the
                * config_byte_counter
                */
                config_byte_counter <= 0;
                // Signal that a new configuration is available
                new_config_available <= 1;
            end else begin
                // A complete byte has been received
                config_byte_counter <= config_byte_counter + 1;
            end
        end else begin
            new_config_available <= 0;
        end
    end
end

/*
 * Process for the transmission part of the spi slave
 * The Hall module sends rotation data to this module, then
 * it needs to send it back through spi_miso to the SBC.
 */

always_ff @(posedge spi_clk or negedge nrst) begin
    if (~nrst) begin
        transmit_register <= DEFAULT_CONFIG_DATA;
        transmission_step <= NO_TRANSMISSION;
    end else begin
        if (~spi_ss) begin
            if (shift_counter == 7) begin
                if ({receive_register[6:0], spi_mosi} == ROTATION_COMMAND) begin
                    transmit_register <= rotation_data[7:0];
                    transmission_step <= FIRST_BYTE;
                end else if (transmission_step == 1) begin
                    transmit_register <= rotation_data[15:8];
                    transmission_step <= SECOND_BYTE;
                end else if (transmission_step == 2) begin
                    transmission_step <= NO_TRANSMISSION;
                end
            end else begin
                transmit_register <= {transmit_register[6:0],1'b1};
            end
        end else begin
            transmit_register[7] <= 1;
        end
    end
end

endmodule
