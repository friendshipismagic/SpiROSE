// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

module EP3C40
(
// {ALTERA_ARGS_BEGIN} DO NOT REMOVE THIS LINE!

	GPIO1,
	GPIO2,
	GPIO3,
	GPIO4,
	GPIO5,
	GPIO6,
	GPIO7,
	GPIO8,
	GPIO9,
	GPIO10,
	GPIO11,
	GPIO12,
	GPIO13,
	GPIO14,
	GPIO15,
	GPIO16,
	GPIO17,
	GPIO18,
	GPIO19,
	GPIO20,
	GPIO21,
	GPIO22,
	GPIO23,
	GPIO24,
	GPIO25,
	GPIO26,
	GPIO27,
	GPIO28,
	GPIO29,
	GPIO30,
	GPIO31,
	GPIO32,
	GPIO33,
	GPIO34,
	GPIO35,
	GPIO36,
	GPIO37,
	GPIO38,
	GPIO39,
	GPIO40,
	GPIO41,
	GPIO42,
	GPIO43,
	GPIO44,
	GPIO45,
	GPIO46,
	GPIO47,
	GPIO48,
	GPIO49,
	GPIO50,
	GPIO51,
	GPIO52,
	GPIO53,
	GPIO54,
	GPIO55,
	GPIO56,
	GPIO57,
	GPIO58,
	GPIO59,
	GPIO60,
	GPIO61,
	GPIO62,
	GPIO63,
	GPIO64,
	GPIO65,
	GPIO66,
	GPIO67,
	GPIO68,
	GPIO69,
	GPIO70,
	GPIO71,
	GPIO72,
	GPIO73,
	GPIO74,
	GPIO75,
	GPIO76,
	GPIO77,
	GPIO78,
	GPIO79,
	GPIO80,
	GPIO81,
	GPIO82,
	GPIO83,
	GPIO84,
	GPIO85,
	GPIO86,
	GPIO87,
	GPIO88,
	GPIO89,
	GPIO90,
	GPIO91,
	GPIO92,
	GPIO93,
	GPIO94,
	GPIO95,
	GPIO96,
	GPIO97,
	GPIO98,
	GPIO99,
	GPIO100,
	GPIO101,
	GPIO102,
	GPIO103
// {ALTERA_ARGS_END} DO NOT REMOVE THIS LINE!

);

// {ALTERA_IO_BEGIN} DO NOT REMOVE THIS LINE!
inout			GPIO1;
inout			GPIO2;
input			GPIO3;
inout			GPIO4;
input			GPIO5;
inout			GPIO6;
inout			GPIO7;
inout			GPIO8;
inout			GPIO9;
inout			GPIO10;
inout			GPIO11;
inout			GPIO12;
inout			GPIO13;
inout			GPIO14;
inout			GPIO15;
inout			GPIO16;
inout			GPIO17;
inout			GPIO18;
inout			GPIO19;
inout			GPIO20;
inout			GPIO21;
inout			GPIO22;
inout			GPIO23;
inout			GPIO24;
inout			GPIO25;
inout			GPIO26;
inout			GPIO27;
inout			GPIO28;
inout			GPIO29;
inout			GPIO30;
inout			GPIO31;
inout			GPIO32;
inout			GPIO33;
inout			GPIO34;
inout			GPIO35;
inout			GPIO36;
inout			GPIO37;
inout			GPIO38;
inout			GPIO39;
inout			GPIO40;
inout			GPIO41;
inout			GPIO42;
inout			GPIO43;
inout			GPIO44;
inout			GPIO45;
inout			GPIO46;
inout			GPIO47;
inout			GPIO48;
inout			GPIO49;
inout			GPIO50;
inout			GPIO51;
inout			GPIO52;
inout			GPIO53;
inout			GPIO54;
inout			GPIO55;
inout			GPIO56;
inout			GPIO57;
inout			GPIO58;
inout			GPIO59;
inout			GPIO60;
inout			GPIO61;
inout			GPIO62;
inout			GPIO63;
inout			GPIO64;
inout			GPIO65;
inout			GPIO66;
inout			GPIO67;
inout			GPIO68;
inout			GPIO69;
inout			GPIO70;
inout			GPIO71;
inout			GPIO72;
inout			GPIO73;
inout			GPIO74;
inout			GPIO75;
inout			GPIO76;
inout			GPIO77;
inout			GPIO78;
inout			GPIO79;
inout			GPIO80;
inout			GPIO81;
inout			GPIO82;
inout			GPIO83;
inout			GPIO84;
inout			GPIO85;
inout			GPIO86;
inout			GPIO87;
inout			GPIO88;
inout			GPIO89;
inout			GPIO90;
inout			GPIO91;
inout			GPIO92;
inout			GPIO93;
inout			GPIO94;
inout			GPIO95;
inout			GPIO96;
inout			GPIO97;
inout			GPIO98;
inout			GPIO99;
inout			GPIO100;
inout			GPIO101;
inout			GPIO102;
inout			GPIO103;

// {ALTERA_IO_END} DO NOT REMOVE THIS LINE!
// {ALTERA_MODULE_BEGIN} DO NOT REMOVE THIS LINE!
// {ALTERA_MODULE_END} DO NOT REMOVE THIS LINE!
endmodule




