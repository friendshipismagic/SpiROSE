/*
 * The SPI is used as an interface between the SOM and
 * the FPGA in order to (from the point of view of the FPGA):
 *   - Receive a new configuration for the drivers
 *   - Transmit rotation information given by the Hall effect
 *   sensors to the SBC
 */

module spi_decoder(
    input  nrst,
    input  clk,

    input  valid,
    input  [55:0] cmd_read,
    output [47:0] cmd_write,

    // Data generated by the Hall sensor module
    input [15:0] rotation_data,

    output new_config_available,
    output rgb_enable
);

localparam CONFIG_COMMAND = 'hBF;
localparam ROTATION_COMMAND = 'h4C;
localparam DISABLE_RGB_COMMAND = 'hD0;
localparam ENABLE_RGB_COMMAND = 'hE0;
localparam DEFAULT_CONFIG_DATA = 'hFF;

`include "drivers_conf.sv"

always_ff @(posedge clk or negedge nrst)
    if (~nrst) begin
        new_config_available <= 0;
        configuration <= serialized_conf;
        rgb_enable <= 0;
    end else begin
        new_config_available <= '0;
        if (valid) begin
            if (cmd_read[55:48] == CONFIG_COMMAND) begin
                configuration <= cmd_read[47:0];
                new_config_available <= '1;
            end else if (cmd_read[7:0] == ENABLE_RGB_COMMAND) begin
                rgb_enable <= '1;
            end else if (cmd_read[7:0] == DISABLE_RGB_COMMAND) begin
                rgb_enable <= '0;
            end
        end
    end

endmodule
